--After Unfolding and pipelining
LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use WORK.fir_package.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;

library std;
use std.textio.all;

entity FIR is
  PORT(DIN  : IN signed(nb-1 downto 0);
	    DIN1 : IN signed(nb-1 downto 0);
		 DIN2 : IN signed(nb-1 downto 0);
		 H0 : in signed (nb-1 downto 0);
		 H1 : in signed (nb-1 downto 0);
		 H2 : in signed (nb-1 downto 0);
		 H3 : in signed (nb-1 downto 0);
		 H4 : in signed (nb-1 downto 0);
		 H5 : in signed (nb-1 downto 0);
		 H6 : in signed (nb-1 downto 0);
		 H7 : in signed (nb-1 downto 0);
		 H8 : in signed (nb-1 downto 0);
		 H9 : in signed (nb-1 downto 0);
		 H10 : in signed (nb-1 downto 0);
       VIN : IN std_logic;
       RST_n : IN std_logic;
       CLK : IN std_logic;
       DOUT  : OUT signed(nb-1 downto 0);
		 DOUT1 : OUT signed(nb-1 downto 0);
		 DOUT2 : OUT signed(nb-1 downto 0);
       VOUT : OUT std_logic );
end FIR; 
architecture BEHAVIOR of FIR is

component REG is
	Port (REG_IN    :	In	signed(nb_opt-1 downto 0);
	      REG_EN    :	In	std_logic;
	      REG_CLK   :	In	std_logic;
         REG_RESET :	In	std_logic;
         REG_OUT   : Out signed(nb_opt-1 downto 0));
end component;
component mult_add is
  PORT(M0 : in signed (nb_opt-1 downto 0);
       M1 : in signed (nb_opt-1 downto 0);
		 M2 : in signed (nb_opt-1 downto 0);
		 M3 : in signed (nb_opt-1 downto 0);
		 M4 : in signed (nb_opt-1 downto 0);
		 M5 : in signed (nb_opt-1 downto 0);
		 M6 : in signed (nb_opt-1 downto 0);
		 M7 : in signed (nb_opt-1 downto 0);
		 M8 : in signed (nb_opt-1 downto 0);
		 M9 : in signed (nb_opt-1 downto 0);
		 M10 :in signed (nb_opt-1 downto 0);
		 
		 H0 : in signed (nb_opt-1 downto 0);
		 H1 : in signed (nb_opt-1 downto 0);
		 H2 : in signed (nb_opt-1 downto 0);
		 H3 : in signed (nb_opt-1 downto 0);
		 H4 : in signed (nb_opt-1 downto 0);
		 H5 : in signed (nb_opt-1 downto 0);
		 H6 : in signed (nb_opt-1 downto 0);
		 H7 : in signed (nb_opt-1 downto 0);
		 H8 : in signed (nb_opt-1 downto 0);
		 H9 : in signed (nb_opt-1 downto 0);
		 H10: in signed (nb_opt-1 downto 0);
       
		 VIN_ma : IN std_logic;
       RST_n_ma : IN std_logic;
       CLK_ma : IN std_logic;
       YOUT  : OUT signed(2*nb_opt-1 downto 0));
end component; 

type sig_vector is array (N downto 0) of signed(nb_opt-1 downto 0);
type regsig_vector is array (13 downto 0) of signed (nb_opt-1 downto 0);
signal b_vect   : sig_vector := (others =>(others =>'0'));
signal x_in, x_in1, x_in2 : regsig_vector;-- := (others =>(others =>'0'));
signal y_out, y_out1, y_out2 : signed(2*nb_opt-1 downto 0);
begin
  b_vect(0) <= H0( (nb-1) downto (nb-nb_opt) ); --Consider high nb_opt bits
  b_vect(1) <= H1( (nb-1) downto (nb-nb_opt) );
  b_vect(2) <= H2( (nb-1) downto (nb-nb_opt) );
  b_vect(3) <= H3( (nb-1) downto (nb-nb_opt) );
  b_vect(4) <= H4( (nb-1) downto (nb-nb_opt) );
  b_vect(5) <= H5( (nb-1) downto (nb-nb_opt) );
  b_vect(6) <= H6( (nb-1) downto (nb-nb_opt) );
  b_vect(7) <= H7( (nb-1) downto (nb-nb_opt) );
  b_vect(8) <= H8( (nb-1) downto (nb-nb_opt) );
  b_vect(9) <= H9( (nb-1) downto (nb-nb_opt) );
  b_vect(10)<= H10((nb-1) downto (nb-nb_opt) );


  process(DIN,DIN1,DIN2)
  begin 
    if (VIN = '1') then 
		VOUT <= '1'; --Dout is ready		
        x_in(0) <= DIN( (nb-1) downto (nb-nb_opt) );
        x_in1(0) <= DIN1( (nb-1) downto (nb-nb_opt) );
        x_in2(0) <= DIN2( (nb-1) downto (nb-nb_opt) );
	 else
	   VOUT <= '0';--Dout is not ready
	 end if;
  end process;

--Perform delayed branch
  FF_loop: for i in 0 to 12 generate
     FF_0_i : REG port map(REG_IN => x_in(i) , REG_EN => VIN, REG_CLK => CLK, REG_RESET => RST_n, REG_OUT => x_in(i+1) );
	 FF_1_i : REG port map(REG_IN => x_in1(i), REG_EN => VIN, REG_CLK => CLK, REG_RESET => RST_n, REG_OUT => x_in1(i+1));
	 FF_2_i : REG port map(REG_IN => x_in2(i), REG_EN => VIN, REG_CLK => CLK, REG_RESET => RST_n, REG_OUT => x_in2(i+1));
  end generate;
---------------------------------------------------------------------------------------------------  
--For pipelining

--First branch
MUL_ADD0 : mult_add port map(M0 => x_in(0), M1 => x_in2(1), M2 => x_in1(2), M3 => x_in(3), M4 => x_in2(5), M5 => x_in1(6), 
                    M6 => x_in(7), M7 => x_in2(9), M8 => x_in1(10), M9 => x_in(11), M10 => x_in2(13),
						  H0 => b_vect(0), H1 => b_vect(1), H2 => b_vect(2), H3 => b_vect(3), H4 => b_vect(4), H5 => b_vect(5), 
						  H6 => b_vect(6), H7 => b_vect(7), H8 => b_vect(8), H9 => b_vect(9), H10 => b_vect(10), 
						  VIN_ma => VIN, RST_n_ma => RST_n, CLK_ma => CLK, YOUT => y_out);   
--Second branch
  MUL_ADD1 : mult_add port map(M0 => x_in1(0), M1 => x_in(0), M2 => x_in2(2), M3 => x_in1(3), M4 => x_in(4), M5 => x_in2(6), 
                    M6 => x_in1(7), M7 => x_in(8), M8 => x_in2(10), M9 => x_in1(11), M10 => x_in(12),
						  H0 => b_vect(0), H1 => b_vect(1), H2 => b_vect(2), H3 => b_vect(3), H4 => b_vect(4), H5 => b_vect(5), 
						  H6 => b_vect(6), H7 => b_vect(7), H8 => b_vect(8), H9 => b_vect(9), H10 => b_vect(10), 

                               						  VIN_ma => VIN, RST_n_ma => RST_n, CLK_ma => CLK, YOUT => y_out1);   
--Third branch
  MUL_ADD2 : mult_add port map(M0 => x_in2(0), M1 => x_in1(0), M2 => x_in(1), M3 => x_in2(3), M4 => x_in1(4), M5 => x_in(5), 
                    M6 => x_in2(7), M7 => x_in1(8), M8 => x_in(9), M9 => x_in2(11), M10 => x_in1(12),
						  H0 => b_vect(0), H1 => b_vect(1), H2 => b_vect(2), H3 => b_vect(3), H4 => b_vect(4), H5 => b_vect(5), 
						  H6 => b_vect(6), H7 => b_vect(7), H8 => b_vect(8), H9 => b_vect(9), H10 => b_vect(10), 
						  VIN_ma => VIN, RST_n_ma => RST_n, CLK_ma => CLK, YOUT => y_out2);   

-------------------------------------------------------------------------------------------------------------
--No pipeline
--First branch
--  MUL_ADD0 : mult_add port map(M0 => x_in(0), M1 => x_in2(1), M2 => x_in1(1), M3 => x_in(1), M4 => x_in2(2), M5 => x_in1(2), 
--                    M6 => x_in(2), M7 => x_in2(3), M8 => x_in1(3), M9 => x_in(3), M10 => x_in2(4),
--						  H0 => b_vect(0), H1 => b_vect(1), H2 => b_vect(2), H3 => b_vect(3), H4 => b_vect(4), H5 => b_vect(5), 
--						  H6 => b_vect(6), H7 => b_vect(7), H8 => b_vect(8), H9 => b_vect(9), H10 => b_vect(10), 
--						  VIN_ma => VIN, RST_n_ma => RST_n, CLK_ma => CLK, YOUT => y_out);   
--Second branch
--  MUL_ADD1 : mult_add port map(M0 => x_in1(0), M1 => x_in(0), M2 => x_in2(1), M3 => x_in1(1), M4 => x_in(1), M5 => x_in2(2), 
--                    M6 => x_in1(2), M7 => x_in(2), M8 => x_in2(3), M9 => x_in1(3), M10 => x_in(3),
--						  H0 => b_vect(0), H1 => b_vect(1), H2 => b_vect(2), H3 => b_vect(3), H4 => b_vect(4), H5 => b_vect(5), 
--						  H6 => b_vect(6), H7 => b_vect(7), H8 => b_vect(8), H9 => b_vect(9), H10 => b_vect(10), 
--						  VIN_ma => VIN, RST_n_ma => RST_n, CLK_ma => CLK, YOUT => y_out1);   
--Third branch
--  MUL_ADD2 : mult_add port map(M0 => x_in2(0), M1 => x_in1(0), M2 => x_in(0), M3 => x_in2(1), M4 => x_in1(1), M5 => x_in(1), 
--                    M6 => x_in2(2), M7 => x_in1(2), M8 => x_in(2), M9 => x_in2(3), M10 => x_in1(3),
--						  H0 => b_vect(0), H1 => b_vect(1), H2 => b_vect(2), H3 => b_vect(3), H4 => b_vect(4), H5 => b_vect(5), 
--						  H6 => b_vect(6), H7 => b_vect(7), H8 => b_vect(8), H9 => b_vect(9), H10 => b_vect(10), 
--						  VIN_ma => VIN, RST_n_ma => RST_n, CLK_ma => CLK, YOUT => y_out2);   

  DOUT  <= y_out( nb-1 downto 0) sll (nb-nb_opt);
  DOUT1 <= y_out1(nb-1 downto 0) sll (nb-nb_opt);
  DOUT2 <= y_out2(nb-1 downto 0) sll (nb-nb_opt);

end BEHAVIOR;
