LIBRARY ieee;
use ieee.std_logic_vector.all;
use ieee.numeric_std.all;

PACKAGE fir_package is
  
  constant nb : integer := 8;
  constant N : integer := 10;

END PACKAGE;
